module scoreDisplay(clk, reset, score, hexsign, hexscore);
	
	input logic clk, reset;
	input logic signed [6:0] score;
	output logic [6:0] hexsign, hexscore;
	
	
	
endmodule 